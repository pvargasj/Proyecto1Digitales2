`include "phy_tx_cond.v" 		

module phy_cond(
    input [7:0] data_in_0_c,
    input [7:0] data_in_1_c,
    input valid_in_0_c,
    input valid_in_1_c,
    input clk_f,
    input clk_2f,
    input clk_8f,
    input reset,
);


endmodule